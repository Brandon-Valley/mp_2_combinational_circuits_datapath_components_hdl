// -- python C:\Users\Brandon\Documents\Personal_Projects\my_utils\modelsim_utils\auto_run.py -d run_cmd__NAND4_v.do

module NOT1_v
  (input i_a,
   output o_f);
   
  assign o_f = ~i_a;
  
endmodule







