// -- python C:\Users\Brandon\Documents\Personal_Projects\my_utils\modelsim_utils\auto_run.py -d run_cmd__NAND4_v.do

module NAND2_v
  (input i_a, i_b,
   output o_f);
   
  assign o_f = ~(i_a & i_b);
  
endmodule







