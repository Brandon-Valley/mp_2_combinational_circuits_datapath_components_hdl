


module OR2_v
  (input i_a, i_b,
   output o_f);
   
  assign o_f = i_a | i_b;
  
  endmodule